`include "defines.v"
//现场可编程IO整列
module fpioa (
    input wire clk,
    input wire rst_n,

    input wire[7:0] waddr_i,
    input wire[`MemBus] data_i,
    input wire[3:0] sel_i,
    input wire we_i,
    input wire[7:0] raddr_i,
    input wire rd_i,
    output reg[`MemBus] data_o,

	input wire [31:0]gpio_oe,//输出使能
	input wire [31:0]gpio_out,//输出数据
    output wire [31:0]gpio_in,//输入数据

    inout wire [31:0] fpioa//处理器IO接口
);
/*------------------------------
 * 线网配置方案
 * 32个FPIOA与256个外设端口互联，形成现场可编程IO整列
 * 
 * 1. 输入数据: fpioa -> 外设
 * 32个FPIOA通过选择器，全部相或，输出至唯一外设端口
 * 
 * 2. 输出数据: 外设 -> fpioa; 输出使能: 外设 -> fpioa
 * 256个外设端口，通过256选1多路选择器，输出至唯一FPIOA端口
 * 
 * 特性：每个FPIOA端口，对应唯一外设端口
 * 每个外设端口，可以同时连接多个FPIOA端口
*/

/*------------------------------
 * 外设端口布局
 * 最大支持256个外设端口，外设端口0恒为空端口
 * 端口布局由 [Number/编号] [Function/功能] [描述] 构成，布局列表如下：
 * | Number   | Function        | 描述                      
 * |----------|-----------------|------------------------------------
 * | 0        | Null            | FPIOA端口默认状态，高阻，输入输出无效
 * | 1        | SPI0_SCK        | 
 * | 2        | SPI0_MOSI       | 
 * | 3        | SPI0_MISO       | 
 * | 4        | SPI0_CS         | 
 * | 5        |                 | 
 * | 6        |                 | 
 * | 7        |                 | 
 * | 8        |                 | 
 * | 9        |                 | 
 * | 10       |                 | 
 * | 11       |                 | 
 * | 12       |                 | 
 * | 13       |                 | 
 * | 14       |                 | 
 * | 15       |                 | 
 * | 16       |                 | 
 * | 17       |                 | 
 * | 18       |                 | 
 * | 19       |                 | 
 * | 20       |                 | 
 * | 21       |                 | 
 * | 22       |                 | 
 * | 23       |                 | 
 * | 24       |                 | 
 * | 25       |                 | 
 * | 26       |                 | 
 * | 27       |                 | 
 * | 28       |                 | 
 * | 29       |                 | 
 * | 30       |                 | 
 * | 31       |                 | 
 * | 32       |                 | 
 * | 33       |                 | 
 * | 34       |                 | 
 * | 35       |                 | 
 * | 36       |                 | 
 * | 37       |                 | 
 * | 38       |                 | 
 * | 39       |                 | 
 * | 40       |                 | 
 * | 41       |                 | 
 * | 42       |                 | 
 * | 43       |                 | 
 * | 44       |                 | 
 * | 45       |                 | 
 * | 46       |                 | 
 * | 47       |                 | 
 * | 48       |                 | 
 * | 49       |                 | 
 * | 50       |                 | 
 * | 51       |                 | 
 * | 52       |                 | 
 * | 53       |                 | 
 * | 54       |                 | 
 * | 55       |                 | 
 * | 56       |                 | 
 * | 57       |                 | 
 * | 58       |                 | 
 * | 59       |                 | 
 * | 60       |                 | 
 * | 61       |                 | 
 * | 62       |                 | 
 * | 63       |                 | 
 * | 64       |                 | 
 * | 65       |                 | 
 * | 66       |                 | 
 * | 67       |                 | 
 * | 68       |                 | 
 * | 69       |                 | 
 * | 70       |                 | 
 * | 71       |                 | 
 * | 72       |                 | 
 * | 73       |                 | 
 * | 74       |                 | 
 * | 75       |                 | 
 * | 76       |                 | 
 * | 77       |                 | 
 * | 78       |                 | 
 * | 79       |                 | 
 * | 80       |                 | 
 * | 81       |                 | 
 * | 82       |                 | 
 * | 83       |                 | 
 * | 84       |                 | 
 * | 85       |                 | 
 * | 86       |                 | 
 * | 87       |                 | 
 * | 88       |                 | 
 * | 89       |                 | 
 * | 90       |                 | 
 * | 91       |                 | 
 * | 92       |                 | 
 * | 93       |                 | 
 * | 94       |                 | 
 * | 95       |                 | 
 * | 96       |                 | 
 * | 97       |                 | 
 * | 98       |                 | 
 * | 99       |                 | 
 * | 100      |                 | 
 * | 101      |                 | 
 * | 102      |                 | 
 * | 103      |                 | 
 * | 104      |                 | 
 * | 105      |                 | 
 * | 106      |                 | 
 * | 107      |                 | 
 * | 108      |                 | 
 * | 109      |                 | 
 * | 110      |                 | 
 * | 111      |                 | 
 * | 112      |                 | 
 * | 113      |                 | 
 * | 114      |                 | 
 * | 115      |                 | 
 * | 116      |                 | 
 * | 117      |                 | 
 * | 118      |                 | 
 * | 119      |                 | 
 * | 120      |                 | 
 * | 121      |                 | 
 * | 122      |                 | 
 * | 123      |                 | 
 * | 124      |                 | 
 * | 125      |                 | 
 * | 126      |                 | 
 * | 127      |                 | 
 * | 128      |                 | 
 * | 129      |                 | 
 * | 130      |                 | 
 * | 131      |                 | 
 * | 132      |                 | 
 * | 133      |                 | 
 * | 134      |                 | 
 * | 135      |                 | 
 * | 136      |                 | 
 * | 137      |                 | 
 * | 138      |                 | 
 * | 139      |                 | 
 * | 140      |                 | 
 * | 141      |                 | 
 * | 142      |                 | 
 * | 143      |                 | 
 * | 144      |                 | 
 * | 145      |                 | 
 * | 146      |                 | 
 * | 147      |                 | 
 * | 148      |                 | 
 * | 149      |                 | 
 * | 150      |                 | 
 * | 151      |                 | 
 * | 152      |                 | 
 * | 153      |                 | 
 * | 154      |                 | 
 * | 155      |                 | 
 * | 156      |                 | 
 * | 157      |                 | 
 * | 158      |                 | 
 * | 159      |                 | 
 * | 160      |                 | 
 * | 161      |                 | 
 * | 162      |                 | 
 * | 163      |                 | 
 * | 164      |                 | 
 * | 165      |                 | 
 * | 166      |                 | 
 * | 167      |                 | 
 * | 168      |                 | 
 * | 169      |                 | 
 * | 170      |                 | 
 * | 171      |                 | 
 * | 172      |                 | 
 * | 173      |                 | 
 * | 174      |                 | 
 * | 175      |                 | 
 * | 176      |                 | 
 * | 177      |                 | 
 * | 178      |                 | 
 * | 179      |                 | 
 * | 180      |                 | 
 * | 181      |                 | 
 * | 182      |                 | 
 * | 183      |                 | 
 * | 184      |                 | 
 * | 185      |                 | 
 * | 186      |                 | 
 * | 187      |                 | 
 * | 188      |                 | 
 * | 189      |                 | 
 * | 190      |                 | 
 * | 191      |                 | 
 * | 192      |                 | 
 * | 193      |                 | 
 * | 194      |                 | 
 * | 195      |                 | 
 * | 196      |                 | 
 * | 197      |                 | 
 * | 198      |                 | 
 * | 199      |                 | 
 * | 200      |                 | 
 * | 201      |                 | 
 * | 202      |                 | 
 * | 203      |                 | 
 * | 204      |                 | 
 * | 205      |                 | 
 * | 206      |                 | 
 * | 207      |                 | 
 * | 208      |                 | 
 * | 209      |                 | 
 * | 210      |                 | 
 * | 211      |                 | 
 * | 212      |                 | 
 * | 213      |                 | 
 * | 214      |                 | 
 * | 215      |                 | 
 * | 216      |                 | 
 * | 217      |                 | 
 * | 218      |                 | 
 * | 219      |                 | 
 * | 220      |                 | 
 * | 221      |                 | 
 * | 222      |                 | 
 * | 223      |                 | 
 * | 224      |                 | 
 * | 225      |                 | 
 * | 226      |                 | 
 * | 227      |                 | 
 * | 228      |                 | 
 * | 229      |                 | 
 * | 230      |                 | 
 * | 231      |                 | 
 * | 232      |                 | 
 * | 233      |                 | 
 * | 234      |                 | 
 * | 235      |                 | 
 * | 236      |                 | 
 * | 237      |                 | 
 * | 238      |                 | 
 * | 239      |                 | 
 * | 240      |                 | 
 * | 241      |                 | 
 * | 242      |                 | 
 * | 243      |                 | 
 * | 244      |                 | 
 * | 245      |                 | 
 * | 246      |                 | 
 * | 247      |                 | 
 * | 248      |                 | 
 * | 249      |                 | 
 * | 250      |                 | 
 * | 251      |                 | 
 * | 252      |                 | 
 * | 253      |                 | 
 * | 254      |                 | 
 * | 255      |                 | 
 * |----------|-----------------|------------------------------------
*/
assign gpio_in = fpioa;
//GPIO中断
genvar i;
for (i = 0; i<32; i=i+1) begin
    assign fpioa[i] = gpio_oe[i] ? gpio_out[i] : 1'bz;
end

wire [255:0]fpioa_sw[0:31];//位宽256，对应256个外设。深度32，对应32个IO口

// 寄存器(偏移)地址
localparam GPIO_DIN = 8'h0;//输入数据
localparam GPIO_OPT = 8'h4;//输出数据
localparam GPIO_OEC = 8'h8;//输出使能
localparam GPIO_TAI = 8'hc;//外部中断控制
/*


// 输入数据，只读
// [31:0]对应GPIO0-31的当前的高低电平
reg [31:0] gpio_din;

// 输出数据，读写
// [31:0]对应GPIO0-31的输出值
reg [31:0] gpio_opt;

// 输出使能，读写
// [31:0]对应GPIO0-31的输出使能状态
reg [31:0] gpio_oec;

// 输出数据，读写
// GPIO0-15的外部中断使能与控制
// [x*2]:  GPIOx中断使能
// [x*2+1]:GPIOx中断为 1:高电平, 2:低电平触发
reg [31:0] gpio_tai;

// 总线接口 写
always @ (posedge clk or negedge rst_n) begin
    if (~rst_n) begin
        gpio_opt <= 32'h0;
        gpio_oec <= 32'h0;
		gpio_tai <= 32'h0;
    end else begin
        if (we_i == 1'b1) begin
            case (waddr_i[3:0])
                GPIO_DIN: ;
				GPIO_OPT: gpio_opt <= data_i;
				GPIO_OEC: gpio_oec <= data_i;
				GPIO_TAI: gpio_tai <= data_i;
                default: ;
            endcase
        end 
		else begin

        end
    end
end

// 总线接口 读
always @ (posedge clk) begin
    if (rd_i == 1'b1) begin
        case (raddr_i[3:0])
                GPIO_DIN: data_o <= gpio_din;
				GPIO_OPT: data_o <= gpio_opt;
				GPIO_OEC: data_o <= gpio_oec;
				GPIO_TAI: data_o <= gpio_tai;
            default: begin
                data_o <= 32'h0;
            end
        endcase
    end
    else begin
        data_o <= data_o;
    end
end

*/


endmodule