module bootrom (
	input clk,    // Clock

	
);

endmodule