module bootrom (
	input wire clk,    // Clock
	input wire [9:0] addr,
	input wire en,
	output [31:0] dout
);

endmodule